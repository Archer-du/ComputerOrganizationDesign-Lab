module SEG_REG(
);
endmodule